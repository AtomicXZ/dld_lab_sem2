module myAnd(input1, input2, op);
  input input1, input2;
  output op;
  and(op, input1, input2);
endmodule