module myNand(input1, input2, op);
	input input1, input2;
	output op;
	nand(op, input1, input2);
endmodule