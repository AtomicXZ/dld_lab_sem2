module myOr(input1, input2, op);
	input input1, input2;
	output op;
	or(op, input1, input2);
endmodule